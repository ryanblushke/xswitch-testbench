/*
  Ryan Blushke, ryb861, 11177824
  CME 435 - 01, Fall Term 2019
  Project, December 5, 2019
*/
program automatic testbench(downstream.driver dstreams[4], upstream.monitor ustreams[4]);
  initial begin
    $display("******************* Start of testcase ****************");
  end

  final
    $display("******************* End of testcase ****************");
endprogram
